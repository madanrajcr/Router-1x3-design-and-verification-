

`define RAM_WIDTH 64
`define ADDR_SIZE 12

typedef enum bit { BAD_XTN,GOOD_XTN}addr_t; 
